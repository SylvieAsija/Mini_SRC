`timescale 1ns/1ns

module boothMultiplier_tb;

reg [31:0] a, b;
wire [63:0] c;

boothMultiplier multiply(a,b,c);

initial
	begin
		a = 2;
		b = 2;
		#10
		a = 0;
		b = 0;
		
	end
	
endmodule