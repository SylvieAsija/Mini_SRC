module incPC(input wire [31:0] a, output wire [31:0] result);

    assign result = a + 1;
    
endmodule