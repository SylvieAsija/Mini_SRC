module bitRecodingMultiplier(input [31:0] in_M, in_Q, output [31:0] out_product)

    

endmodule