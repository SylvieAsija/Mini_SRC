//module ALU(input [31:0] controlSignal, input YMuxIn, BusIn, output [31:0] out)

    

//endmodule