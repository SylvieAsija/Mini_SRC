module Encoder(output reg [4:0] out, input [31:0] data);
	always@(*)
	begin
		if(data == 32'b00000000000000000000000000000001) out = 0; else
		if(data == 32'b00000000000000000000000000000010) out = 1; else
		if(data == 32'b00000000000000000000000000000100) out = 2; else
		if(data == 32'b00000000000000000000000000001000) out = 3; else
		if(data == 32'b00000000000000000000000000010000) out = 4; else
		if(data == 32'b00000000000000000000000000100000) out = 5; else
		if(data == 32'b00000000000000000000000001000000) out = 6; else
		if(data == 32'b00000000000000000000000010000000) out = 7; else
		if(data == 32'b00000000000000000000000100000000) out = 8; else
		if(data == 32'b00000000000000000000001000000000) out = 9; else
		if(data == 32'b00000000000000000000010000000000) out = 10; else
		if(data == 32'b00000000000000000000100000000000) out = 11; else
		if(data == 32'b00000000000000000001000000000000) out = 12; else
		if(data == 32'b00000000000000000010000000000000) out = 13; else
		if(data == 32'b00000000000000000100000000000000) out = 14; else
		if(data == 32'b00000000000000001000000000000000) out = 15; else
		if(data == 32'b00000000000000010000000000000000) out = 16; else
		if(data == 32'b00000000000000100000000000000000) out = 17; else
		if(data == 32'b00000000000001000000000000000000) out = 18; else
		if(data == 32'b00000000000010000000000000000000) out = 19; else
		if(data == 32'b00000000000100000000000000000000) out = 20; else
		if(data == 32'b00000000001000000000000000000000) out = 21; else
		if(data == 32'b00000000010000000000000000000000) out = 22; else
		if(data == 32'b00000000100000000000000000000000) out = 23; else
		if(data == 32'b00000001000000000000000000000000) out = 24; else
		if(data == 32'b00000010000000000000000000000000) out = 25; else
		if(data == 32'b00000100000000000000000000000000) out = 26; else
		if(data == 32'b00001000000000000000000000000000) out = 27; else
		if(data == 32'b00010000000000000000000000000000) out = 28; else
		if(data == 32'b00100000000000000000000000000000) out = 29; else
		if(data == 32'b01000000000000000000000000000000) out = 30; else
		if(data == 32'b10000000000000000000000000000000) out = 31; else out = 5'bx;
		
	end
endmodule
