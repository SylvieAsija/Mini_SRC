module memoryDataRegister(input [31:0] BusMuxOut, Mdatain, output [31:0] out, input read, clear, clock, MDRin)
    

endmodule