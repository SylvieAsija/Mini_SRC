module memoryDataRegister(input [31:0] BusMuxOut, Mdatain, output [31:0] BusMuxIn-MDR, memChip, input read, clear, clock, MDRin)


endmodule